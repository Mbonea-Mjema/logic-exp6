library verilog;
use verilog.vl_types.all;
entity Vend_FSM_vlg_vec_tst is
end Vend_FSM_vlg_vec_tst;
